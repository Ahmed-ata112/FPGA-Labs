��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��$�����Q�-E�zW�l5n$�0��4WO�G&z��|��T�<��r��Xz�q�*���*i�В-L_O�B��pL����V����d��Gc]%��u���c��D����G��G��F����������zAO49��4��r�~2��u`���Q�9�h�����tdFM)f���a'(�*�S]Oޫ,UL�.	�3v����=�V�g1�efjl@@@�7<�<m���JЅ}^e�m��9�"�j�(��'�y0hT�T�B�qfz9߆��'�
�x�p-�7zK�ёt��*��|\��	 <���z��OF�`�����ׯ�������9C��@��f�+�#&��\7|��K|�g�Mh莸?>��~�BM�D���'�g/s�a���z$5[ZՍ���]�6�m���'��u��t�I\36��������x���<m���z�]�3�_?���yC�0~�k�y1��=T��qд��]@5U������Ų���2Տ�\��{���J�����)"���`�vD���q�og~U���5V���'�B2CP���X���1�^�ir��qR)�̛���������Q}@l�t���&]0�W*-`b�g�D	��16��0�pGe�~��N/�������|�f��7mk��l��c�q���vYфrǔ��7�Z�f>B��@��q.؃�A�/�L�y��׭���(+�Z��8�nv��dX@�^�w�}=�v�uJ0}�r�����#��0mQ��Կ�i�4����/�|G�b�@���7���@\��� �m���T�bR�\�]=V�i�ʓh�.Ƃn�Ơ[�=�r�?!���V��6)K`C�З����"e[ꥠ�TK�.��Q�"Gx�
�ì�=T��m��<$��p�b� �+4���+X"�H!7����p��MpYL�(�7���Q�ϵm�Wd�T/��Lm��Hj��������&�T^�UH_IG��h���Ҏ�r
=�J�S7��[�; �r~��-��@�%!-���*!P#��Z��~��e�#!+B��3�;3�����Q��l��B}�I�حs�"F|�������Wv�XE[�9�CJT�K�~�>��\�θ �G�
��?9*t�>c5ꐏ��]<Y
�3��󌥍�G��G\���wDWܪA��0��ݲ6XM&P�3�g{/sJ�R�x���X%��s����F}����6z�K��"11�ޚ���և<Ro���
�f�
7�%c?I`$q�}�#�C�Pm��]�6��ݔ�Y���4�P������]�Ӯ{]_�)�����w
���v���4|}f�H��b�{����qr��.E��bG��&�zm(���pK0�X��I��-�i��"o�G2����D$]&m[Y��O�Q�T��4WUT��t������4�W_��z����wM����ӟ�(�I֜��q���%�a��#�i^r��q�'���}����0ر,���Skr $d�j�5��q�pJ��G�(�����R�<�Z��<��l*M�S����&�8�U�{x�&��'�+]���t�CH&�!�?\Hy���֊8G�Uk`D���;����8U��"��-��{B���#��{|��	� �s���N���], k�'q��,�9u�t�1ˣ܅h/0�l���2��B�rO��HO�=���F6+�\�-�7�8� ��~0����QM�-z���Z��-�<�[%���"��'��C�G���JLLb%ߕ� �ծ�?|���oɶWE�N�QE�\`�3��ӊI���2EgN*BY!��/ ũُ��QG�i���p���'"Ğ��3�L9���!�S�O�^�|ƆC h�6�k���L�'%�����F������h�ҫ7��D��|cT�{p���ڝ2��3l�����BP��c��[tUt�q��1���R'V���@8���X�;x�e�����M$�Y"s|mW1�5�D�A�P��Kj� �������7і��o?)�%f�i#^;~\�T�#$��}�^�P F�~�����˩�@����kD}ܚu�z�l#�]�
��ܾ�%!��i\���$n� ��&�Q��2W���=I9���.С�6��n�Bz�F�2�<�9_l
�!P����τʢħ�)H�`���&�\�%y;��J#d�K �}池7`�(#"�mV�3��X�F4[�rަ�M������좲���<��/%�f��j-Vi�D)�EEu��7�ec�[B��mY|�~�W��� +,'���vÆ����/I
�4����J{ :�5�b�r�Fb��rG����YqO2�����!Ƶ�s��������ì�_��	\5qB��mcpyV���{5YwƉ�f>�=fԖ7��6�y1�*�-��%�ѥ�r{�0D���*'FZ002���v�;ד*{e������6&(�M��	\���G�(��\�6Ű�_P5�"���$c��q�%f9�sP����w뚭�bH��Z�*1�
�C�2�8	,w�`�K��\7y��,��w)�a��m	om�ڦ;�!��g�S���TR�]�K�`
��,�חo0T��2{#�v]e|�<%d��Fl�
}����(r�%�=�?�t�Y��9��O_�3��r����߳&��>
h��H�ϩ��,B$n�d0�������Q���z�vbה�&��i~F����7�	~���|y�����N=۳�4�_G��B��k�߫cD��n�ᛜ�B���+��bzg�; ��)�R�s��7���١"�S7�/Z:���䈮c"��$��V^S����Hi�����z]��� �#��úY����WCȓ^޿UWbDNk\G�Q2=�unChص^֤*��t�}�̋�-�	��Z+�H,w�������a
T l��U
���� 3��,zVvPBIZ���$Ҝ��r?�&k�޾c�������Di�<C�lq=���T_�P1@��ѦX��I,蘴�������(,��9�]m��x?_i��/l?b ;��>L�y1��{F�����U/U���oӹ��!�C����rEފ�_o�M�	@!oC��^	{u��D�4�S;E^#I�.��n+����y{Z�	�P/��z���R���t;#V56ıt,�5�\B�(�2�����:K����� 2ylX)f����h�Sz��.�jԦ���Z�
O:	�xy�"�kš�K͔sW�yݤu�q�=f��Ez�7�"b�Wz���N��G��]�?tZf~������z�,߁Q�&�7�D�&=X�x��o�����Vw��H�1�����^d}��fr�Aza ("��80l������k�D/���Ø��	������5�ѯ�&ܬHW ���p�vCb���&���ǠWc0����*�4K���<����a�Lħ��C�l�6�@̴�;��p]�(/:�O��o�*;�*Ux���Y�1+؆\"��>��|��G���D�}�?���oW��������{嬣+�� A����3����SBz�Έ}ۊ��
bW�9m���ߙ��WL��j�Z&�ÍkJ��nC*;�}�x��˪�/Bi=t����(����*�s��>�|��Z(h�3���Q�� �g-�دn�%$��6����2�ٹd�)���\{GI_)f�A���+����5�B��Lfj(��՟��:fr��c�O�Q����L|����5�M.�u�1��EOK;�n
,���ڽ�|�Ͽ_[��M#r�f0�Ǡ#��Ϗ�¢���zP��%�M�Dq烷EoF������,���g%��_�@�|�ޛs��*Epˈh���K�V���u�te�CpT*~�t�Pm� k�.,K�p4�:m����*I�O/��8Y�ؘݹ�q������noV�w�KY$?Î���Fy4�',Z�u�pA
,�{���˷K}�b�,Pcnl }��|�D,��L�
��{��Fw�ʋ>����s�v��9�G����Ұ��=m$�X�I]r8a!�_������l2��M�ͧ���������&^�T�ה�sc�Mwa+ `?�^F�B5CU;?����=��= �;��y��!ܿ�yt��=�\�,���E�G?Z�>t�X�(J�1g�!r�ZY��za<f��̬��1H��Ɋej;���A%�����L��BY�(<�c�	L�!�'Z@��#3^%&�b�6�����/�ǀ���x�@�F
�!�#E�������E���sê�*�䓦��J!��妡$�sXU�}d�,I]}a���%�R�5�u�Q#��鼞3O\�/�ncG��h=���]Ac+�0M�6bF2�� �*�'�iɶ�5�r�0)�98P�l%�V��R�g��+\'(M,�Fł5I���^Ta�*�P��'z�M�V�ܬ�rOg��Kɺ_��X5�C�57�VT[����-K��N��E� ]q.���n~Umf��/��H^��/�I�[g[��q�|�&Pv���U11v��;��u����Q�GT�4��%	;{4]����݇&��z�ޱ����CX�v\���RA�]��sЬ��xF	���i:���>��{�R�bh�~$5��
Y���k㎃G��6�i,�d�r���_�o�*��g`��Z3(6�~ҵ��-���yL���+iUd���q���f٘
/���/!Yn�=gT�K���o�m��U�3��a횃�'������!��| 0�_��,qm�*�����qX6�:q/Ĵd�M�Z�h�T������,4/#bpotŷ�ԋ�����/����2i�sFr���z;簹U�j����k[J�j��o���8����HR,�~�]�ۇr�J lna�H<:����@@M� H�D��l�¼�J]����(���bX��ˍ%k����a�j�Q��Z���Y�Y],}�Ts���L���v��Z��Q\��c,�t���,��t8n�m���A"��OoKL*v�}�zբ�sW9���g���y�4�&B��`��5%mf5ٖMn]�� tW%j#WE�c�Эism���wE� O0�Âo%X}�TI�W+���ڐ��쫯���b���N��n����g0��+,!��n��TsJb|���v��~���������uU�N���=�V�L�J頠3в5�J˴M�p��zfϾ%���k{k��|�H��m�u ���i�l0��V��k��>�K��%@>��`)��7ݛk�
xo�6�c~��Z������Ժ�[��O��Q��	\�'
�Vg�2�o%�G+. RG�A˥�q�7Z�K7������Rp�[���lWs�Pj�_�K5��ڋD�ۻ.LMW���2�h��s2N�/R�������j@�-_��6�10I	K L����W@�����۰Q���@��M/9��P�2c�2�B�Q�I?\���v}�n��bc��M�Q�>Q��jQՃ9�*��S-I�I�_���v�섰^�F��y&0�t��Q�ð�P+����W�ևcH�A���r�����K�S��I>؍�ԛ�l<}����;6��x�����EneQ�V��|�f�!�QQ���'Y�EQ$F&sZ����-��s'��08�(Q�X��.& �,��Lg@Q��m�x⪝��=k������s�K�l���lhD�����[�6>�ʎA��NfC�)�d�RI�L���0�$��1�^����+b#��u��>&��=>���H^���ԫ�H7;ֿ�>�y8R�́��QQb�--�%�UԱ,�$�ս&b�R����p7}.
, �<$���o�:w�r|��8Հ\h_�8���@���:-�L���b��B�Z^�$���*�4�.��}�"[��{
��&!z��(h�6�F��DA�#'���1����35��|�z_�[�l��Air"�*��2�{�7Н��VN?��+�4��9�4?XQ���S�wdr;G��|��KI���4~�
T��a^���&�7
F�0=䦪�W�a��v�kvA�b��޵���g��[#.�ݹ��!VN���*t���y0����#^;��ɷ�����a�L!�wO��[]-��U�0�p�3*7�����$4���%(lZrwfn��#9�9h×������n�A݋���=H�픝Dˆ�̛Kh{�?纙 ڛ�j.,xjB�C��<��_f���~�&�"�2��R���t�_^=�*ɖ�~�{$�}�c�e�R�`���.(�Zy����<����e0��8	�'���U��iv?V{���V_��M�q��2�N�i�(q���8�	a4�5�c�j+N�w��DE��1�����ߔ�Hȋ3�ʚ��x3%X1D\�%��d�%���fy���۔������=|k��|����2����\��S6c���a��Mm����J
����`�^0_��prZ�����#�Y��hN	�����H|��X�F ��݉�^�lRk^���%rU�D��6�t=~H&��������~djs��MF���^�.��ۉ�t�xAL&��~~���� ��5'f�J��ѽ:�nj����_��P�R��N��և �2\��.#y��WF5}�_�>FK��~ ��w�`��߆iT���1Aɪ#��=���Տ3X�L?ܶR�X�]P>�X���KH	e��ox$�M��m�{=����Wơ�i��yߊ����,���C�O�(�@#�0Y�E`�<B?��_Qeq]t��Uv
��R�-���. ���C��P�-if^Ų���ŉE'\M߱�x�Oy���>�]PG���t_Z��b-
���9N�$�ܾ�e>��<��4ǯD�zn��U���򚗼!9���=��F�a��*�~�Ji��^����/����DqDt�c�b�?�|���U��fpf�`1�����"�J] �̚'�U覢n�/?�PR����lҙ�U��/������LKP��5*�9�&��W#�o�����3��zn����q�g ���E����6 �,i'D���siH����KY�h���e�X��b���ıA9�%�9|����<C_�����i�To��	V�F6�%p��!����ڣx��R㵅����SX݋�����$bZ汝�s�j�������*�f3Z��5\9?���K���\/� �za9b�$q�~����#��+�AQd.����.�T��̵����q��׆ȥ!�:},��GY��t��=�wVg����qK4�m�6N�V��Z݁V�jk0h��q�f�e˸Cnw�_���c��4ߑ���١���)O�r�qs��`c���z�=!�sF}��o
<V�M���?�Fg)�	cÀv@�U���?���&�\A�ӯ�Ge]�\��\����+htb�˂Eh�+²2��ّ�%jI�r�/�4ݓlK��v�>��`�j�j��۵�C�;vh!6�Az�4�	kk�c�RG�`)I��U�bm��k�Sh�6X0��MHr�-& Ǒ2�Q�u\�N^��3�o$�%wI٣�r���\�ʑkP�]�)|��t��{c19е�R��iCm����Ȧ��~�+XSV�.3��9h�j��^����l�	+�v�D�t2������z�[�P����.�i��nj�D:~�O��P�װ�uS��S��5ؿ��R�!Ԑ����2?�EnkyX4:ޣ4#`���G ��d�u��kSIS���1�?�V};�j'�Ͷb�Y����S��QUF���Q���?�� ��׿b��ZԶ�Y5��y�����9��,0�IC�f�u��D[�>$�����col[HO�
vpj���F��'��Y[�B]���]�V����ݪ��q���v�8�T6�r���F�σ��fֆ�X&-p8z��]S�@��}�<���,��EhU�o��*�;�5I����2�ӨP������/�$��8�׀�[6��[ng�	�\��x[���5m�\wY����zW��&Q�vn�)�=����5�G��cÔR�����[b}�uQ�-�T`�\����8����B�Y�4�C��y��S<α�%�7��Է݀�0��Ed�J�VgW�d���;L��RDdʊ,:�(h����K��ƥ�DO��p����������^�u��K
����K�K��?��)D~���6T�&V�-�]_-�V�F宵?kױ!��c�aE��O'5P���g/T�t�p�����bQ(�dӜ��x�ʜ�.4=j��i���:����/7=��չ��5UGD����)6}��%��]eC�����U*A�!gZồk��:�t�ޕ�*҆�PCx�O�#�!����x�+#�G�Y�
�)Ȇ�,M��H-R".�8��q"poG����$��im��]���㿑����x���Rf�/�wШ�˩�%�p�p@��a�_�K�n#�h�"��m�]�K@~p)���[�ކ0��i���,S�	nw����dy��
�D�=_�����b�w\e12	G/��o�!����	Z�2}�OH>%��IꍠN����ׇ���h�) �z�o&Ā�A`{�Z�(\N��A+R��`u�o��J����17'��薘%͜�*T��[˻��ۻ��0����-|$��V1��Z��+㞜u�M�@d��#MG7���T\笜�U��)��|P����5�l�N5�����e�x{�vR�_�s'���J��H��tN��}>Qi���Xg#�Q�ٺ�p�2�q����?	bdZ�q\��D���k�
����i�~c#Mp�L��l|k#�̋ �B�P-�-wL����R�ʠA Ԝ�Yj@축j�E}˞���2H�М��P8�nC9�/���~����DK�|�3B� A\ʧ�|]����t{~����7Q`\�EOw#9��V��|N��O������Xt���lǠ�l���$Wd�s�5�g^���	}���
�J_SJ���Q�a�.�Ǣ*0S6ݚ�W�z�em��P��'���X2��XPZbSMb����o�B4
j���(�:`��&�4���4�/jH͎�`��Ո}~��J\)�C��3j��+ߠX���;ށ�qk8&��MP�����q�]�M�;'��Vg#���n�hf/_3�>W��Z#�.p V������,�S�����sw;�q�!�&ΙGe�8�4��@5�� �{m�p���n���dMBH��V�$4��
v䀺�- ��s�9j� K�O`��}����I�?|1��Νok�S|�By֟�U�/�K[}n� � �\����*�&u�|�p�9�0�Gs"�ULq���",�?0��c�_}��̷Р�NJ��0_և�T`������
�	5�%�!�2a]a������9o?�֤�G�@ˏ)�_�`:�*����*ƹ�M����a�`<��2����W�s[*��j$�dX��G|d.�:��/?�O�!�v�6�^+��Aə��ա��7�RpnuGP�'�Q�g|hƷ�0ZD�SZ����4��Yu����֯֦�HL*�)����8A���Q%BG���)�	P�%��<\M�"(zԓ��V�419~^9y2�y6�<�5!~�3�ɂ����kU��O��/M. ��&���!�z=Z!��!|B-ktR��v2��}Bx��KO��b�/��'QG�c�� \IW8�b����`4����?R�G�x�[P�doT�1����z^ß�;�`��	����+�p�%�������R
o��&A�a���b�L�f�Q�j]�k��G�K�ժ���G���  �V��d;�S���S�՛XMF
g��*�M��mՙ�hv��i��pR4��wF��I{_�	O)&uyX��BBl�4y�{/0���.(�A�D ���
�#�6Տ�?~��Yf�HI�
����T�/���TaQ��'�|�s�u(�\��W=|p��?Tag]��w�ȭwX[D����ǕS���&?v��x�-��&C�����b(qJ�п���D,������v���0o�="������D���=}��%����>�	PntT��?���;��K[ʸl��ִ�@ƴ*ȸ�k�yGѠ[���rV�Ak⨏=�%E��k�K ~�����N�<*���lf�ş87��r�<��-.?�=I�{4���Sƍ���9׀<�60�7Q,��Fu�@tD�Rǘ����tm?�A�F�8T��t�;���|*5T}W���68��W����x�摞��˨bs8�S�A	l�mc\��z�$*�r�O	$�Lu:2T/����f�2p򿫯��tg�{�+������i������D��dw)*�����.�.�M�T�X)�7�xA#��ZF0��ȴ����Q0�E���� ��b]�U7^i��K���RH79��v�\�e�l�zBH�V�%�R"Si߶�Y	(Pa!�^�����pA?|a�|�S��c%t���`W�"sW���r�y���}2�*$$l1-��-�X܇��}�ATz�i��P����, ܖ�ib�?5�;5^)~(ar��g����@c�~5�
�?�s��C���] �׊�Ci����
�-���&���1K�R���;�گ�� �-��+,�����%޴A�i{����@r,8��f���',�yܚ|��R�o��`�_��X[g����aU��_�/�O�j��G�euû�+݂�%~y4��O��6{�*A]�0f��|* ������[�R�#馡\.5��*7�a�)�c+*c[W�`N����~3�Ԋ3�u�i���^�����%�Ea7|�2�ȧ�`ZDכ�>��-�_�\�c_;��5-�UY���m%�h.ݳ5Ms[0�eu$�y��2�R/�)��>����D�ό>y`��i�p��D��rsR�s��@�vz�~��@��Yi�D�c���ҟUs��N�ܵh8!d��6��â|����Q�e31֨�t>ϵ��)&��Iə��,J�/���f�t!�a�D�#�Qj�]�"���J�CV��cw�y?\����l� �S�6�e�b���v��Lt�{�aLw^����e�W�:�M��dK"��.V�_���\!�y.��|sr�����o	4Pq>Td �c=�ҏ��u����)��M]�f s2Eάs����L!ʗ�z�o��Zy�WT�ɕR���֊��U�w�"��[���_|^{�3L'��z��˽�* �M�'%g�fe���ƀs�O�]o�ir�5C��h=��T��m���w.�^�Uȿ�%ᇰ=`�譓�@V%�9�Su[��y��3; V%���%��$5����PO�\o�R��(j�����<d
�e�6��Q0����q,u�0f���^��`8�B/�jb�\}��'-�O�_5�I���jN�&ط��)C���u��{��,�C*_��T�춺������6|��5ֽ��f���%�q���){[tE�w�+���O��dDVp��5�*j�f����i�ŝ\!���kz��en�h�C�|l�ŏ�V��ݬ��d������uHG��R�~X��ZK6جѾ��ȓҰH�{j�j��d�P�_������Mn��V�?Jr��K�[Zm!�1�S����2s�˖A��_��{l1�-�K%��A9��L��4���V�a�\�I"����$gTF��{��آgP7�i缆}*�tqQTs;H9ը�8J���2RQF����6�dT�>��D�@��u͡�6ڷ4�{br.��0�-&y%v��b�ʦ(�K����F�n#uT�Ԏ��^��<k8\�1�7��a��N���_����>}Kqtۇʧ�`
/d���	M8f��F�S��.B���qf�� �c��@�|���i�~���"G@� ��ԩ�/�[��fw�pΧ��bQ{iz�&�<����*�y�F�}'��}�dVnT���{���bF��ϰ����,y�~3V����t,�X�^�ȯ�B-0�V�b"��=@�	��g�:�(ORWm����:���R�{[N 6z��>��D�+�#�է�c�Ln��>3C�� ]C3~�=\��Y���F��Z�w 
DG�&�Aj������